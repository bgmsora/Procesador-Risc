LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ExtensorSigno IS

	PORT (

		ENTRADA : IN STD_LOGIC_VECTOR(11 DOWNTO 0);

		SALIDA : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)

	);

END ExtensorSigno;

ARCHITECTURE Arquitectura OF ExtensorSigno IS

	SIGNAL MSB : STD_LOGIC;

BEGIN

	MSB <= ENTRADA(11);

	SALIDA <= MSB & MSB & MSB & MSB & ENTRADA;

END Arquitectura;